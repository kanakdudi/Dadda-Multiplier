module stage1_16to13 (
    input  [15:0] PP16_1,
    input  [15:0] PP16_2,
    input  [15:0] PP16_3,
    input  [15:0] PP16_4,
    input  [15:0] PP16_5,
    input  [15:0] PP16_6,
    input  [15:0] PP16_7,
    input  [15:0] PP16_8,
    input  [15:0] PP16_9,
    input  [15:0] PP16_10,
    input  [15:0] PP16_11,
    input  [15:0] PP16_12,
    input  [15:0] PP16_13,
    input  [15:0] PP16_14,
    input  [15:0] PP16_15,
    input  [15:0] PP16_16,
    output [30:0] PP13_1,
    output [29:1] PP13_2,
    output [28:2] PP13_3,
    output [27:3] PP13_4,
    output [26:4] PP13_5,
    output [25:5] PP13_6,
    output [24:6] PP13_7,
    output [23:7] PP13_8,
    output [22:8] PP13_9,
    output [21:9] PP13_10,
    output [20:10] PP13_11,
    output [19:11] PP13_12,
    output [19:12] PP13_13
);
    wire S13_ha, C13_ha;
    wire S14_fa1, C14_fa1, S14_ha1, C14_ha1;
    wire S15_fa1, C15_fa1, S15_fa2, C15_fa2, S15_ha1, C15_ha1;
    wire S16_fa1, C16_fa1, S16_fa2, C16_fa2, S16_fa3, C16_fa3;
    wire S17_fa1, C17_fa1, S17_fa2, C17_fa2;
    wire S18_fa1, C18_fa1;

    
    // 13th column
    HA ha13_1 ( .A(PP16_1[13]), .B(PP16_2[12]), .Sum(S13_ha), .Cout(C13_ha));

    // 14th column
    FA fa14_1 ( .A(PP16_1[14]), .B(PP16_2[13]), .Cin(PP16_3[12]), .Sum(S14_fa1), .Cout(C14_fa1));
    HA ha14_1 ( .A(PP16_5[10]), .B(PP16_4[11]), .Sum(S14_ha1), .Cout(C14_ha1));

    // 15th column
    FA fa15_1 ( .A(PP16_1[15]), .B(PP16_2[14]), .Cin(PP16_3[13]), .Sum(S15_fa1), .Cout(C15_fa1));
    FA fa15_2 ( .A(PP16_4[12]), .B(PP16_5[11]), .Cin(PP16_6[10]), .Sum(S15_fa2), .Cout(C15_fa2));
    HA ha15_1 ( .A(PP16_7[9]), .B(PP16_8[8]), .Sum(S15_ha1), .Cout(C15_ha1));

    // 16th column

    /* 
    FA fa16_1 ( .A(PP16_2[15]), .B(PP16_3[14]), .Cin(PP16_4[13]), .Sum(S16_fa1), .Cout(C16_fa1));
    FA fa16_2 ( .A(PP16_5[12]), .B(PP16_6[11]), .Cin(PP16_7[10]), .Sum(S16_fa2), .Cout(C16_fa2));
    FA fa16_3 ( .A(PP16_8[9]), .B(PP16_9[8]), .Cin(PP16_10[7]), .Sum(S16_fa3), .Cout(C16_fa3));
     */

    FA fa16_1 ( .A(PP16_2[15]), .B(PP16_3[14]), .Cin(1'b1), .Sum(S16_fa1), .Cout(C16_fa1));
    FA fa16_2 ( .A(PP16_4[13]), .B(PP16_5[12]), .Cin(PP16_6[11]), .Sum(S16_fa2), .Cout(C16_fa2));
    FA fa16_3 ( .A(PP16_7[10]), .B(PP16_9[8]), .Cin(PP16_8[9]), .Sum(S16_fa3), .Cout(C16_fa3));

    // 17th column
    FA fa17_1 ( .A(PP16_3[15]), .B(PP16_4[14]), .Cin(PP16_5[13]), .Sum(S17_fa1), .Cout(C17_fa1));
    FA fa17_2 ( .A(PP16_6[12]), .B(PP16_7[11]), .Cin(PP16_8[10]), .Sum(S17_fa2), .Cout(C17_fa2)); 

    // 18th column
    FA fa18_1 ( .A(PP16_4[15]), .B(PP16_5[14]), .Cin(PP16_6[13]), .Sum(S18_fa1), .Cout(C18_fa1));  


    // Assign outputs
    assign PP13_1[30:0] = {PP16_16[15], PP16_15[15], PP16_14[15], PP16_13[15], PP16_12[15], PP16_11[15], PP16_10[15], PP16_9[15], PP16_8[15], PP16_7[15], PP16_6[15], C18_fa1, C17_fa1, C16_fa1, C15_fa1, C14_fa1, C13_ha, S13_ha, PP16_1[12:0]}; 
    assign PP13_2[29:1] = {PP16_16[14], PP16_15[14], PP16_14[14], PP16_13[14], PP16_12[14], PP16_11[14], PP16_10[14], PP16_9[14], PP16_8[14], PP16_7[14], PP16_5[15], C17_fa2, C16_fa2, C15_fa2, C14_ha1, S14_fa1, PP16_3[11], PP16_2[11:0]};
    assign PP13_3[28:2] = {PP16_16[13], PP16_15[13], PP16_14[13], PP16_13[13], PP16_12[13], PP16_11[13], PP16_10[13], PP16_9[13], PP16_8[13], PP16_6[14], S18_fa1, C16_fa3, C15_ha1, S15_fa1, S14_ha1, PP16_4[10], PP16_3[10:0]};
    assign PP13_4[27:3] = {PP16_16[12], PP16_15[12], PP16_14[12], PP16_13[12], PP16_12[12], PP16_11[12], PP16_10[12], PP16_9[12], PP16_7[13], PP16_7[12], S17_fa1, S16_fa1, S15_fa2, PP16_6[9], PP16_5[9], PP16_4[9:0]};
    assign PP13_5[26:4] = {PP16_16[11], PP16_15[11], PP16_14[11], PP16_13[11], PP16_12[11], PP16_11[11], PP16_10[11], PP16_8[12], PP16_8[11], S17_fa2, S16_fa2, S15_ha1, PP16_7[8], PP16_6[8], PP16_5[8:0]};
    assign PP13_6[25:5] = {PP16_16[10], PP16_15[10], PP16_14[10], PP16_13[10], PP16_12[10], PP16_11[10], PP16_9[11], PP16_9[10], PP16_9[9], S16_fa3, PP16_9[7], PP16_8[7], PP16_7[7], PP16_6[7:0]};
    assign PP13_7[24:6] = {PP16_16[9], PP16_15[9], PP16_14[9], PP16_13[9], PP16_12[9], PP16_10[10], PP16_10[9], PP16_10[8], PP16_10[7], PP16_10[6], PP16_9[6], PP16_8[6], PP16_7[6:0]};
    assign PP13_8[23:7] = {PP16_16[8], PP16_15[8], PP16_14[8], PP16_13[8], PP16_11[9], PP16_11[8], PP16_11[7], PP16_11[6], PP16_11[5], PP16_10[5], PP16_9[5], PP16_8[5:0]};
    assign PP13_9[22:8] = {PP16_16[7], PP16_15[7], PP16_14[7], PP16_12[8], PP16_12[7], PP16_12[6], PP16_12[5], PP16_12[4], PP16_11[4], PP16_10[4], PP16_9[4:0]};
    assign PP13_10[21:9] = {PP16_16[6], PP16_15[6], PP16_13[7], PP16_13[6], PP16_13[5], PP16_13[4], PP16_13[3], PP16_12[3], PP16_11[3], PP16_10[3:0]};
    assign PP13_11[20:10] = {PP16_16[5], PP16_14[6], PP16_14[5], PP16_14[4], PP16_14[3], PP16_14[2], PP16_13[2], PP16_12[2], PP16_11[2:0]};
    assign PP13_12[19:11] = {PP16_15[5], PP16_15[4], PP16_15[3], PP16_15[2], PP16_15[1], PP16_14[1], PP16_13[1], PP16_12[1:0]};
    assign PP13_13[19:12] = {PP16_16[4], PP16_16[3], PP16_16[2], PP16_16[1], PP16_16[0], PP16_15[0], PP16_14[0], PP16_13[0]};

 
 endmodule